// megafunction wizard: %Shift register (RAM-based)%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTSHIFT_TAPS 

// ============================================================
// File Name: count_sr.v
// Megafunction Name(s):
// 			ALTSHIFT_TAPS
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 23.1std.0 Build 991 11/28/2023 SC Lite Edition
// ************************************************************

//Copyright (C) 2023  Intel Corporation. All rights reserved.
//Your use of Intel Corporation's design tools, logic functions 
//and other software and tools, and any partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Intel Program License 
//Subscription Agreement, the Intel Quartus Prime License Agreement,
//the Intel FPGA IP License Agreement, or other applicable license
//agreement, including, without limitation, that your use is for
//the sole purpose of programming logic devices manufactured by
//Intel and sold by Intel or its authorized distributors.  Please
//refer to the applicable agreement for further details, at
//https://fpgasoftware.intel.com/eula.

module count_sr (
	clock,
	shiftin,
	shiftout,
	taps);

	input	  clock;
	input	[20:0]  shiftin;
	output	[20:0]  shiftout;
	output	[20:0]  taps;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: ACLR NUMERIC "0"
// Retrieval info: PRIVATE: CLKEN NUMERIC "0"
// Retrieval info: PRIVATE: GROUP_TAPS NUMERIC "0"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: PRIVATE: NUMBER_OF_TAPS NUMERIC "1"
// Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "0"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: TAP_DISTANCE NUMERIC "6"
// Retrieval info: PRIVATE: WIDTH NUMERIC "21"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: CONSTANT: LPM_HINT STRING "RAM_BLOCK_TYPE=MLAB"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altshift_taps"
// Retrieval info: CONSTANT: NUMBER_OF_TAPS NUMERIC "1"
// Retrieval info: CONSTANT: TAP_DISTANCE NUMERIC "6"
// Retrieval info: CONSTANT: WIDTH NUMERIC "21"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
// Retrieval info: USED_PORT: shiftin 0 0 21 0 INPUT NODEFVAL "shiftin[20..0]"
// Retrieval info: USED_PORT: shiftout 0 0 21 0 OUTPUT NODEFVAL "shiftout[20..0]"
// Retrieval info: USED_PORT: taps 0 0 21 0 OUTPUT NODEFVAL "taps[20..0]"
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @shiftin 0 0 21 0 shiftin 0 0 21 0
// Retrieval info: CONNECT: shiftout 0 0 21 0 @shiftout 0 0 21 0
// Retrieval info: CONNECT: taps 0 0 21 0 @taps 0 0 21 0
// Retrieval info: GEN_FILE: TYPE_NORMAL count_sr.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL count_sr.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL count_sr.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL count_sr.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL count_sr_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL count_sr_bb.v TRUE
// Retrieval info: LIB_FILE: altera_mf
